// soc.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module soc (
		input  wire        clk_clk,            //          clk.clk
		input  wire [31:0] hps_f2h_irq0_irq,   // hps_f2h_irq0.irq
		input  wire [10:0] mem1_s1_address,    //      mem1_s1.address
		input  wire        mem1_s1_clken,      //             .clken
		input  wire        mem1_s1_chipselect, //             .chipselect
		input  wire        mem1_s1_write,      //             .write
		output wire [15:0] mem1_s1_readdata,   //             .readdata
		input  wire [15:0] mem1_s1_writedata,  //             .writedata
		input  wire [1:0]  mem1_s1_byteenable, //             .byteenable
		input  wire [10:0] mem2_s1_address,    //      mem2_s1.address
		input  wire        mem2_s1_clken,      //             .clken
		input  wire        mem2_s1_chipselect, //             .chipselect
		input  wire        mem2_s1_write,      //             .write
		output wire [15:0] mem2_s1_readdata,   //             .readdata
		input  wire [15:0] mem2_s1_writedata,  //             .writedata
		input  wire [1:0]  mem2_s1_byteenable, //             .byteenable
		output wire [14:0] memory_mem_a,       //       memory.mem_a
		output wire [2:0]  memory_mem_ba,      //             .mem_ba
		output wire        memory_mem_ck,      //             .mem_ck
		output wire        memory_mem_ck_n,    //             .mem_ck_n
		output wire        memory_mem_cke,     //             .mem_cke
		output wire        memory_mem_cs_n,    //             .mem_cs_n
		output wire        memory_mem_ras_n,   //             .mem_ras_n
		output wire        memory_mem_cas_n,   //             .mem_cas_n
		output wire        memory_mem_we_n,    //             .mem_we_n
		output wire        memory_mem_reset_n, //             .mem_reset_n
		inout  wire [31:0] memory_mem_dq,      //             .mem_dq
		inout  wire [3:0]  memory_mem_dqs,     //             .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,   //             .mem_dqs_n
		output wire        memory_mem_odt,     //             .mem_odt
		output wire [3:0]  memory_mem_dm,      //             .mem_dm
		input  wire        memory_oct_rzqin,   //             .oct_rzqin
		input  wire        reset_reset_n       //        reset.reset_n
	);

	wire   [1:0] hps_h2f_axi_master_awburst;           // hps:h2f_AWBURST -> mm_interconnect_0:hps_h2f_axi_master_awburst
	wire   [3:0] hps_h2f_axi_master_arlen;             // hps:h2f_ARLEN -> mm_interconnect_0:hps_h2f_axi_master_arlen
	wire   [7:0] hps_h2f_axi_master_wstrb;             // hps:h2f_WSTRB -> mm_interconnect_0:hps_h2f_axi_master_wstrb
	wire         hps_h2f_axi_master_wready;            // mm_interconnect_0:hps_h2f_axi_master_wready -> hps:h2f_WREADY
	wire  [11:0] hps_h2f_axi_master_rid;               // mm_interconnect_0:hps_h2f_axi_master_rid -> hps:h2f_RID
	wire         hps_h2f_axi_master_rready;            // hps:h2f_RREADY -> mm_interconnect_0:hps_h2f_axi_master_rready
	wire   [3:0] hps_h2f_axi_master_awlen;             // hps:h2f_AWLEN -> mm_interconnect_0:hps_h2f_axi_master_awlen
	wire  [11:0] hps_h2f_axi_master_wid;               // hps:h2f_WID -> mm_interconnect_0:hps_h2f_axi_master_wid
	wire   [3:0] hps_h2f_axi_master_arcache;           // hps:h2f_ARCACHE -> mm_interconnect_0:hps_h2f_axi_master_arcache
	wire         hps_h2f_axi_master_wvalid;            // hps:h2f_WVALID -> mm_interconnect_0:hps_h2f_axi_master_wvalid
	wire  [29:0] hps_h2f_axi_master_araddr;            // hps:h2f_ARADDR -> mm_interconnect_0:hps_h2f_axi_master_araddr
	wire   [2:0] hps_h2f_axi_master_arprot;            // hps:h2f_ARPROT -> mm_interconnect_0:hps_h2f_axi_master_arprot
	wire   [2:0] hps_h2f_axi_master_awprot;            // hps:h2f_AWPROT -> mm_interconnect_0:hps_h2f_axi_master_awprot
	wire  [63:0] hps_h2f_axi_master_wdata;             // hps:h2f_WDATA -> mm_interconnect_0:hps_h2f_axi_master_wdata
	wire         hps_h2f_axi_master_arvalid;           // hps:h2f_ARVALID -> mm_interconnect_0:hps_h2f_axi_master_arvalid
	wire   [3:0] hps_h2f_axi_master_awcache;           // hps:h2f_AWCACHE -> mm_interconnect_0:hps_h2f_axi_master_awcache
	wire  [11:0] hps_h2f_axi_master_arid;              // hps:h2f_ARID -> mm_interconnect_0:hps_h2f_axi_master_arid
	wire   [1:0] hps_h2f_axi_master_arlock;            // hps:h2f_ARLOCK -> mm_interconnect_0:hps_h2f_axi_master_arlock
	wire   [1:0] hps_h2f_axi_master_awlock;            // hps:h2f_AWLOCK -> mm_interconnect_0:hps_h2f_axi_master_awlock
	wire  [29:0] hps_h2f_axi_master_awaddr;            // hps:h2f_AWADDR -> mm_interconnect_0:hps_h2f_axi_master_awaddr
	wire   [1:0] hps_h2f_axi_master_bresp;             // mm_interconnect_0:hps_h2f_axi_master_bresp -> hps:h2f_BRESP
	wire         hps_h2f_axi_master_arready;           // mm_interconnect_0:hps_h2f_axi_master_arready -> hps:h2f_ARREADY
	wire  [63:0] hps_h2f_axi_master_rdata;             // mm_interconnect_0:hps_h2f_axi_master_rdata -> hps:h2f_RDATA
	wire         hps_h2f_axi_master_awready;           // mm_interconnect_0:hps_h2f_axi_master_awready -> hps:h2f_AWREADY
	wire   [1:0] hps_h2f_axi_master_arburst;           // hps:h2f_ARBURST -> mm_interconnect_0:hps_h2f_axi_master_arburst
	wire   [2:0] hps_h2f_axi_master_arsize;            // hps:h2f_ARSIZE -> mm_interconnect_0:hps_h2f_axi_master_arsize
	wire         hps_h2f_axi_master_bready;            // hps:h2f_BREADY -> mm_interconnect_0:hps_h2f_axi_master_bready
	wire         hps_h2f_axi_master_rlast;             // mm_interconnect_0:hps_h2f_axi_master_rlast -> hps:h2f_RLAST
	wire         hps_h2f_axi_master_wlast;             // hps:h2f_WLAST -> mm_interconnect_0:hps_h2f_axi_master_wlast
	wire   [1:0] hps_h2f_axi_master_rresp;             // mm_interconnect_0:hps_h2f_axi_master_rresp -> hps:h2f_RRESP
	wire  [11:0] hps_h2f_axi_master_awid;              // hps:h2f_AWID -> mm_interconnect_0:hps_h2f_axi_master_awid
	wire  [11:0] hps_h2f_axi_master_bid;               // mm_interconnect_0:hps_h2f_axi_master_bid -> hps:h2f_BID
	wire         hps_h2f_axi_master_bvalid;            // mm_interconnect_0:hps_h2f_axi_master_bvalid -> hps:h2f_BVALID
	wire   [2:0] hps_h2f_axi_master_awsize;            // hps:h2f_AWSIZE -> mm_interconnect_0:hps_h2f_axi_master_awsize
	wire         hps_h2f_axi_master_awvalid;           // hps:h2f_AWVALID -> mm_interconnect_0:hps_h2f_axi_master_awvalid
	wire         hps_h2f_axi_master_rvalid;            // mm_interconnect_0:hps_h2f_axi_master_rvalid -> hps:h2f_RVALID
	wire         mm_interconnect_0_mem1_s2_chipselect; // mm_interconnect_0:mem1_s2_chipselect -> mem1:chipselect2
	wire  [31:0] mm_interconnect_0_mem1_s2_readdata;   // mem1:readdata2 -> mm_interconnect_0:mem1_s2_readdata
	wire   [9:0] mm_interconnect_0_mem1_s2_address;    // mm_interconnect_0:mem1_s2_address -> mem1:address2
	wire   [3:0] mm_interconnect_0_mem1_s2_byteenable; // mm_interconnect_0:mem1_s2_byteenable -> mem1:byteenable2
	wire         mm_interconnect_0_mem1_s2_write;      // mm_interconnect_0:mem1_s2_write -> mem1:write2
	wire  [31:0] mm_interconnect_0_mem1_s2_writedata;  // mm_interconnect_0:mem1_s2_writedata -> mem1:writedata2
	wire         mm_interconnect_0_mem1_s2_clken;      // mm_interconnect_0:mem1_s2_clken -> mem1:clken2
	wire         mm_interconnect_0_mem2_s2_chipselect; // mm_interconnect_0:mem2_s2_chipselect -> mem2:chipselect2
	wire  [31:0] mm_interconnect_0_mem2_s2_readdata;   // mem2:readdata2 -> mm_interconnect_0:mem2_s2_readdata
	wire   [9:0] mm_interconnect_0_mem2_s2_address;    // mm_interconnect_0:mem2_s2_address -> mem2:address2
	wire   [3:0] mm_interconnect_0_mem2_s2_byteenable; // mm_interconnect_0:mem2_s2_byteenable -> mem2:byteenable2
	wire         mm_interconnect_0_mem2_s2_write;      // mm_interconnect_0:mem2_s2_write -> mem2:write2
	wire  [31:0] mm_interconnect_0_mem2_s2_writedata;  // mm_interconnect_0:mem2_s2_writedata -> mem2:writedata2
	wire         mm_interconnect_0_mem2_s2_clken;      // mm_interconnect_0:mem2_s2_clken -> mem2:clken2
	wire  [31:0] hps_f2h_irq1_irq;                     // irq_mapper:sender_irq -> hps:f2h_irq_p1
	wire         rst_controller_reset_out_reset;       // rst_controller:reset_out -> [mem1:reset, mem2:reset, mm_interconnect_0:mem1_reset1_reset_bridge_in_reset_reset]
	wire         rst_controller_reset_out_reset_req;   // rst_controller:reset_req -> [mem1:reset_req, mem2:reset_req]
	wire         rst_controller_001_reset_out_reset;   // rst_controller_001:reset_out -> mm_interconnect_0:hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	wire         hps_h2f_reset_reset;                  // hps:h2f_rst_n -> rst_controller_001:reset_in0

	soc_hps #(
		.F2S_Width (2),
		.S2F_Width (2)
	) hps (
		.mem_a              (memory_mem_a),               //            memory.mem_a
		.mem_ba             (memory_mem_ba),              //                  .mem_ba
		.mem_ck             (memory_mem_ck),              //                  .mem_ck
		.mem_ck_n           (memory_mem_ck_n),            //                  .mem_ck_n
		.mem_cke            (memory_mem_cke),             //                  .mem_cke
		.mem_cs_n           (memory_mem_cs_n),            //                  .mem_cs_n
		.mem_ras_n          (memory_mem_ras_n),           //                  .mem_ras_n
		.mem_cas_n          (memory_mem_cas_n),           //                  .mem_cas_n
		.mem_we_n           (memory_mem_we_n),            //                  .mem_we_n
		.mem_reset_n        (memory_mem_reset_n),         //                  .mem_reset_n
		.mem_dq             (memory_mem_dq),              //                  .mem_dq
		.mem_dqs            (memory_mem_dqs),             //                  .mem_dqs
		.mem_dqs_n          (memory_mem_dqs_n),           //                  .mem_dqs_n
		.mem_odt            (memory_mem_odt),             //                  .mem_odt
		.mem_dm             (memory_mem_dm),              //                  .mem_dm
		.oct_rzqin          (memory_oct_rzqin),           //                  .oct_rzqin
		.h2f_rst_n          (hps_h2f_reset_reset),        //         h2f_reset.reset_n
		.f2h_sdram0_clk     (clk_clk),                    //  f2h_sdram0_clock.clk
		.f2h_sdram0_ARADDR  (),                           //   f2h_sdram0_data.araddr
		.f2h_sdram0_ARLEN   (),                           //                  .arlen
		.f2h_sdram0_ARID    (),                           //                  .arid
		.f2h_sdram0_ARSIZE  (),                           //                  .arsize
		.f2h_sdram0_ARBURST (),                           //                  .arburst
		.f2h_sdram0_ARLOCK  (),                           //                  .arlock
		.f2h_sdram0_ARPROT  (),                           //                  .arprot
		.f2h_sdram0_ARVALID (),                           //                  .arvalid
		.f2h_sdram0_ARCACHE (),                           //                  .arcache
		.f2h_sdram0_AWADDR  (),                           //                  .awaddr
		.f2h_sdram0_AWLEN   (),                           //                  .awlen
		.f2h_sdram0_AWID    (),                           //                  .awid
		.f2h_sdram0_AWSIZE  (),                           //                  .awsize
		.f2h_sdram0_AWBURST (),                           //                  .awburst
		.f2h_sdram0_AWLOCK  (),                           //                  .awlock
		.f2h_sdram0_AWPROT  (),                           //                  .awprot
		.f2h_sdram0_AWVALID (),                           //                  .awvalid
		.f2h_sdram0_AWCACHE (),                           //                  .awcache
		.f2h_sdram0_BRESP   (),                           //                  .bresp
		.f2h_sdram0_BID     (),                           //                  .bid
		.f2h_sdram0_BVALID  (),                           //                  .bvalid
		.f2h_sdram0_BREADY  (),                           //                  .bready
		.f2h_sdram0_ARREADY (),                           //                  .arready
		.f2h_sdram0_AWREADY (),                           //                  .awready
		.f2h_sdram0_RREADY  (),                           //                  .rready
		.f2h_sdram0_RDATA   (),                           //                  .rdata
		.f2h_sdram0_RRESP   (),                           //                  .rresp
		.f2h_sdram0_RLAST   (),                           //                  .rlast
		.f2h_sdram0_RID     (),                           //                  .rid
		.f2h_sdram0_RVALID  (),                           //                  .rvalid
		.f2h_sdram0_WLAST   (),                           //                  .wlast
		.f2h_sdram0_WVALID  (),                           //                  .wvalid
		.f2h_sdram0_WDATA   (),                           //                  .wdata
		.f2h_sdram0_WSTRB   (),                           //                  .wstrb
		.f2h_sdram0_WREADY  (),                           //                  .wready
		.f2h_sdram0_WID     (),                           //                  .wid
		.h2f_axi_clk        (clk_clk),                    //     h2f_axi_clock.clk
		.h2f_AWID           (hps_h2f_axi_master_awid),    //    h2f_axi_master.awid
		.h2f_AWADDR         (hps_h2f_axi_master_awaddr),  //                  .awaddr
		.h2f_AWLEN          (hps_h2f_axi_master_awlen),   //                  .awlen
		.h2f_AWSIZE         (hps_h2f_axi_master_awsize),  //                  .awsize
		.h2f_AWBURST        (hps_h2f_axi_master_awburst), //                  .awburst
		.h2f_AWLOCK         (hps_h2f_axi_master_awlock),  //                  .awlock
		.h2f_AWCACHE        (hps_h2f_axi_master_awcache), //                  .awcache
		.h2f_AWPROT         (hps_h2f_axi_master_awprot),  //                  .awprot
		.h2f_AWVALID        (hps_h2f_axi_master_awvalid), //                  .awvalid
		.h2f_AWREADY        (hps_h2f_axi_master_awready), //                  .awready
		.h2f_WID            (hps_h2f_axi_master_wid),     //                  .wid
		.h2f_WDATA          (hps_h2f_axi_master_wdata),   //                  .wdata
		.h2f_WSTRB          (hps_h2f_axi_master_wstrb),   //                  .wstrb
		.h2f_WLAST          (hps_h2f_axi_master_wlast),   //                  .wlast
		.h2f_WVALID         (hps_h2f_axi_master_wvalid),  //                  .wvalid
		.h2f_WREADY         (hps_h2f_axi_master_wready),  //                  .wready
		.h2f_BID            (hps_h2f_axi_master_bid),     //                  .bid
		.h2f_BRESP          (hps_h2f_axi_master_bresp),   //                  .bresp
		.h2f_BVALID         (hps_h2f_axi_master_bvalid),  //                  .bvalid
		.h2f_BREADY         (hps_h2f_axi_master_bready),  //                  .bready
		.h2f_ARID           (hps_h2f_axi_master_arid),    //                  .arid
		.h2f_ARADDR         (hps_h2f_axi_master_araddr),  //                  .araddr
		.h2f_ARLEN          (hps_h2f_axi_master_arlen),   //                  .arlen
		.h2f_ARSIZE         (hps_h2f_axi_master_arsize),  //                  .arsize
		.h2f_ARBURST        (hps_h2f_axi_master_arburst), //                  .arburst
		.h2f_ARLOCK         (hps_h2f_axi_master_arlock),  //                  .arlock
		.h2f_ARCACHE        (hps_h2f_axi_master_arcache), //                  .arcache
		.h2f_ARPROT         (hps_h2f_axi_master_arprot),  //                  .arprot
		.h2f_ARVALID        (hps_h2f_axi_master_arvalid), //                  .arvalid
		.h2f_ARREADY        (hps_h2f_axi_master_arready), //                  .arready
		.h2f_RID            (hps_h2f_axi_master_rid),     //                  .rid
		.h2f_RDATA          (hps_h2f_axi_master_rdata),   //                  .rdata
		.h2f_RRESP          (hps_h2f_axi_master_rresp),   //                  .rresp
		.h2f_RLAST          (hps_h2f_axi_master_rlast),   //                  .rlast
		.h2f_RVALID         (hps_h2f_axi_master_rvalid),  //                  .rvalid
		.h2f_RREADY         (hps_h2f_axi_master_rready),  //                  .rready
		.f2h_axi_clk        (clk_clk),                    //     f2h_axi_clock.clk
		.f2h_AWID           (),                           //     f2h_axi_slave.awid
		.f2h_AWADDR         (),                           //                  .awaddr
		.f2h_AWLEN          (),                           //                  .awlen
		.f2h_AWSIZE         (),                           //                  .awsize
		.f2h_AWBURST        (),                           //                  .awburst
		.f2h_AWLOCK         (),                           //                  .awlock
		.f2h_AWCACHE        (),                           //                  .awcache
		.f2h_AWPROT         (),                           //                  .awprot
		.f2h_AWVALID        (),                           //                  .awvalid
		.f2h_AWREADY        (),                           //                  .awready
		.f2h_AWUSER         (),                           //                  .awuser
		.f2h_WID            (),                           //                  .wid
		.f2h_WDATA          (),                           //                  .wdata
		.f2h_WSTRB          (),                           //                  .wstrb
		.f2h_WLAST          (),                           //                  .wlast
		.f2h_WVALID         (),                           //                  .wvalid
		.f2h_WREADY         (),                           //                  .wready
		.f2h_BID            (),                           //                  .bid
		.f2h_BRESP          (),                           //                  .bresp
		.f2h_BVALID         (),                           //                  .bvalid
		.f2h_BREADY         (),                           //                  .bready
		.f2h_ARID           (),                           //                  .arid
		.f2h_ARADDR         (),                           //                  .araddr
		.f2h_ARLEN          (),                           //                  .arlen
		.f2h_ARSIZE         (),                           //                  .arsize
		.f2h_ARBURST        (),                           //                  .arburst
		.f2h_ARLOCK         (),                           //                  .arlock
		.f2h_ARCACHE        (),                           //                  .arcache
		.f2h_ARPROT         (),                           //                  .arprot
		.f2h_ARVALID        (),                           //                  .arvalid
		.f2h_ARREADY        (),                           //                  .arready
		.f2h_ARUSER         (),                           //                  .aruser
		.f2h_RID            (),                           //                  .rid
		.f2h_RDATA          (),                           //                  .rdata
		.f2h_RRESP          (),                           //                  .rresp
		.f2h_RLAST          (),                           //                  .rlast
		.f2h_RVALID         (),                           //                  .rvalid
		.f2h_RREADY         (),                           //                  .rready
		.h2f_lw_axi_clk     (clk_clk),                    //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID        (),                           // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR      (),                           //                  .awaddr
		.h2f_lw_AWLEN       (),                           //                  .awlen
		.h2f_lw_AWSIZE      (),                           //                  .awsize
		.h2f_lw_AWBURST     (),                           //                  .awburst
		.h2f_lw_AWLOCK      (),                           //                  .awlock
		.h2f_lw_AWCACHE     (),                           //                  .awcache
		.h2f_lw_AWPROT      (),                           //                  .awprot
		.h2f_lw_AWVALID     (),                           //                  .awvalid
		.h2f_lw_AWREADY     (),                           //                  .awready
		.h2f_lw_WID         (),                           //                  .wid
		.h2f_lw_WDATA       (),                           //                  .wdata
		.h2f_lw_WSTRB       (),                           //                  .wstrb
		.h2f_lw_WLAST       (),                           //                  .wlast
		.h2f_lw_WVALID      (),                           //                  .wvalid
		.h2f_lw_WREADY      (),                           //                  .wready
		.h2f_lw_BID         (),                           //                  .bid
		.h2f_lw_BRESP       (),                           //                  .bresp
		.h2f_lw_BVALID      (),                           //                  .bvalid
		.h2f_lw_BREADY      (),                           //                  .bready
		.h2f_lw_ARID        (),                           //                  .arid
		.h2f_lw_ARADDR      (),                           //                  .araddr
		.h2f_lw_ARLEN       (),                           //                  .arlen
		.h2f_lw_ARSIZE      (),                           //                  .arsize
		.h2f_lw_ARBURST     (),                           //                  .arburst
		.h2f_lw_ARLOCK      (),                           //                  .arlock
		.h2f_lw_ARCACHE     (),                           //                  .arcache
		.h2f_lw_ARPROT      (),                           //                  .arprot
		.h2f_lw_ARVALID     (),                           //                  .arvalid
		.h2f_lw_ARREADY     (),                           //                  .arready
		.h2f_lw_RID         (),                           //                  .rid
		.h2f_lw_RDATA       (),                           //                  .rdata
		.h2f_lw_RRESP       (),                           //                  .rresp
		.h2f_lw_RLAST       (),                           //                  .rlast
		.h2f_lw_RVALID      (),                           //                  .rvalid
		.h2f_lw_RREADY      (),                           //                  .rready
		.f2h_irq_p0         (hps_f2h_irq0_irq),           //          f2h_irq0.irq
		.f2h_irq_p1         (hps_f2h_irq1_irq)            //          f2h_irq1.irq
	);

	soc_mem1 mem1 (
		.address     (mem1_s1_address),                      //     s1.address
		.clken       (mem1_s1_clken),                        //       .clken
		.chipselect  (mem1_s1_chipselect),                   //       .chipselect
		.write       (mem1_s1_write),                        //       .write
		.readdata    (mem1_s1_readdata),                     //       .readdata
		.writedata   (mem1_s1_writedata),                    //       .writedata
		.byteenable  (mem1_s1_byteenable),                   //       .byteenable
		.address2    (mm_interconnect_0_mem1_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_mem1_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_mem1_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_mem1_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_mem1_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_mem1_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_mem1_s2_byteenable), //       .byteenable
		.clk         (clk_clk),                              //   clk1.clk
		.reset       (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze      (1'b0)                                  // (terminated)
	);

	soc_mem2 mem2 (
		.address     (mem2_s1_address),                      //     s1.address
		.clken       (mem2_s1_clken),                        //       .clken
		.chipselect  (mem2_s1_chipselect),                   //       .chipselect
		.write       (mem2_s1_write),                        //       .write
		.readdata    (mem2_s1_readdata),                     //       .readdata
		.writedata   (mem2_s1_writedata),                    //       .writedata
		.byteenable  (mem2_s1_byteenable),                   //       .byteenable
		.address2    (mm_interconnect_0_mem2_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_mem2_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_mem2_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_mem2_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_mem2_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_mem2_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_mem2_s2_byteenable), //       .byteenable
		.clk         (clk_clk),                              //   clk1.clk
		.reset       (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze      (1'b0)                                  // (terminated)
	);

	soc_mm_interconnect_0 mm_interconnect_0 (
		.hps_h2f_axi_master_awid                                        (hps_h2f_axi_master_awid),              //                                       hps_h2f_axi_master.awid
		.hps_h2f_axi_master_awaddr                                      (hps_h2f_axi_master_awaddr),            //                                                         .awaddr
		.hps_h2f_axi_master_awlen                                       (hps_h2f_axi_master_awlen),             //                                                         .awlen
		.hps_h2f_axi_master_awsize                                      (hps_h2f_axi_master_awsize),            //                                                         .awsize
		.hps_h2f_axi_master_awburst                                     (hps_h2f_axi_master_awburst),           //                                                         .awburst
		.hps_h2f_axi_master_awlock                                      (hps_h2f_axi_master_awlock),            //                                                         .awlock
		.hps_h2f_axi_master_awcache                                     (hps_h2f_axi_master_awcache),           //                                                         .awcache
		.hps_h2f_axi_master_awprot                                      (hps_h2f_axi_master_awprot),            //                                                         .awprot
		.hps_h2f_axi_master_awvalid                                     (hps_h2f_axi_master_awvalid),           //                                                         .awvalid
		.hps_h2f_axi_master_awready                                     (hps_h2f_axi_master_awready),           //                                                         .awready
		.hps_h2f_axi_master_wid                                         (hps_h2f_axi_master_wid),               //                                                         .wid
		.hps_h2f_axi_master_wdata                                       (hps_h2f_axi_master_wdata),             //                                                         .wdata
		.hps_h2f_axi_master_wstrb                                       (hps_h2f_axi_master_wstrb),             //                                                         .wstrb
		.hps_h2f_axi_master_wlast                                       (hps_h2f_axi_master_wlast),             //                                                         .wlast
		.hps_h2f_axi_master_wvalid                                      (hps_h2f_axi_master_wvalid),            //                                                         .wvalid
		.hps_h2f_axi_master_wready                                      (hps_h2f_axi_master_wready),            //                                                         .wready
		.hps_h2f_axi_master_bid                                         (hps_h2f_axi_master_bid),               //                                                         .bid
		.hps_h2f_axi_master_bresp                                       (hps_h2f_axi_master_bresp),             //                                                         .bresp
		.hps_h2f_axi_master_bvalid                                      (hps_h2f_axi_master_bvalid),            //                                                         .bvalid
		.hps_h2f_axi_master_bready                                      (hps_h2f_axi_master_bready),            //                                                         .bready
		.hps_h2f_axi_master_arid                                        (hps_h2f_axi_master_arid),              //                                                         .arid
		.hps_h2f_axi_master_araddr                                      (hps_h2f_axi_master_araddr),            //                                                         .araddr
		.hps_h2f_axi_master_arlen                                       (hps_h2f_axi_master_arlen),             //                                                         .arlen
		.hps_h2f_axi_master_arsize                                      (hps_h2f_axi_master_arsize),            //                                                         .arsize
		.hps_h2f_axi_master_arburst                                     (hps_h2f_axi_master_arburst),           //                                                         .arburst
		.hps_h2f_axi_master_arlock                                      (hps_h2f_axi_master_arlock),            //                                                         .arlock
		.hps_h2f_axi_master_arcache                                     (hps_h2f_axi_master_arcache),           //                                                         .arcache
		.hps_h2f_axi_master_arprot                                      (hps_h2f_axi_master_arprot),            //                                                         .arprot
		.hps_h2f_axi_master_arvalid                                     (hps_h2f_axi_master_arvalid),           //                                                         .arvalid
		.hps_h2f_axi_master_arready                                     (hps_h2f_axi_master_arready),           //                                                         .arready
		.hps_h2f_axi_master_rid                                         (hps_h2f_axi_master_rid),               //                                                         .rid
		.hps_h2f_axi_master_rdata                                       (hps_h2f_axi_master_rdata),             //                                                         .rdata
		.hps_h2f_axi_master_rresp                                       (hps_h2f_axi_master_rresp),             //                                                         .rresp
		.hps_h2f_axi_master_rlast                                       (hps_h2f_axi_master_rlast),             //                                                         .rlast
		.hps_h2f_axi_master_rvalid                                      (hps_h2f_axi_master_rvalid),            //                                                         .rvalid
		.hps_h2f_axi_master_rready                                      (hps_h2f_axi_master_rready),            //                                                         .rready
		.clk_clk_clk                                                    (clk_clk),                              //                                                  clk_clk.clk
		.hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),   // hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.mem1_reset1_reset_bridge_in_reset_reset                        (rst_controller_reset_out_reset),       //                        mem1_reset1_reset_bridge_in_reset.reset
		.mem1_s2_address                                                (mm_interconnect_0_mem1_s2_address),    //                                                  mem1_s2.address
		.mem1_s2_write                                                  (mm_interconnect_0_mem1_s2_write),      //                                                         .write
		.mem1_s2_readdata                                               (mm_interconnect_0_mem1_s2_readdata),   //                                                         .readdata
		.mem1_s2_writedata                                              (mm_interconnect_0_mem1_s2_writedata),  //                                                         .writedata
		.mem1_s2_byteenable                                             (mm_interconnect_0_mem1_s2_byteenable), //                                                         .byteenable
		.mem1_s2_chipselect                                             (mm_interconnect_0_mem1_s2_chipselect), //                                                         .chipselect
		.mem1_s2_clken                                                  (mm_interconnect_0_mem1_s2_clken),      //                                                         .clken
		.mem2_s2_address                                                (mm_interconnect_0_mem2_s2_address),    //                                                  mem2_s2.address
		.mem2_s2_write                                                  (mm_interconnect_0_mem2_s2_write),      //                                                         .write
		.mem2_s2_readdata                                               (mm_interconnect_0_mem2_s2_readdata),   //                                                         .readdata
		.mem2_s2_writedata                                              (mm_interconnect_0_mem2_s2_writedata),  //                                                         .writedata
		.mem2_s2_byteenable                                             (mm_interconnect_0_mem2_s2_byteenable), //                                                         .byteenable
		.mem2_s2_chipselect                                             (mm_interconnect_0_mem2_s2_chipselect), //                                                         .chipselect
		.mem2_s2_clken                                                  (mm_interconnect_0_mem2_s2_clken)       //                                                         .clken
	);

	soc_irq_mapper irq_mapper (
		.clk        (),                 //       clk.clk
		.reset      (),                 // clk_reset.reset
		.sender_irq (hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_h2f_reset_reset),               // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
